module tb_reg;

A_reg (
    .clk,
    .rst_n,
    .a_bus,
    a_cpu,
    a_in,
    a_out
);
endmodule
